//`define USE_LED_FOR_RESET_BLOCK 1
`undef USE_LED_FOR_RESET_BLOCK

//`define USE_LED_FOR_CONFIG_BLOCK 1
`undef USE_LED_FOR_CONFIG_BLOCK

`define USE_LED_FOR_COMM_BLOCK 1
//`undef USE_LED_FOR_COMM_BLOCK



module state_machine(

	// clock and reset
	input 					reset,
	input 					clk, 		// 50 MHz (see https://www.waveshare.com/wiki/OpenEP4CE6-C_User_Manual#Clock_Circuit)
	
	// LEDs
	inout 	reg [3:0]	led,
	
	// ULPI
	input  	wire 			CLKOUT, 	// PIN 50
	input  	wire 			DIR,    	// PIN 52
	input 	wire 			NXT, 		// PIN 54
	output 	wire 			RST,    	// PIN 46	
	output 	reg 			STP, 		// PIN 58	
	inout 	wire [7:0] 	data,
	
	// UART
	output 	wire 			uart_tx_pin, // PIN 
	
	// test
	output 	wire 			TESTPIN

);

	wire 	[7:0] indata;
	reg 	[7:0] outdata;
	
	assign indata = data;
	assign data = DIR ? 8'bz : outdata;
	
	
	
	// when reset is asserted, the phy resets
	reg [31:0] phy_reset_counter;
	reg phy_reset_performed;
	
	reg RST_reg;
	assign RST = RST_reg;

	//reg stp_reg;
	//assign STP = stp_reg;
	
	reg ulpi_register_write_reg;
	
	//reg [3:0] led_reg;
	//assign led = led_reg;
	
	reg [7:0] latched_data_reg;
	
	
	
	//
	// ULPI soft reset logic
	//
	
	// UPLI, Perform RESET
	always @(posedge CLKOUT)
	begin
	
		if (!reset)
		begin
`ifdef USE_LED_FOR_RESET_BLOCK
			led <= ~4'b1110;
`endif

			// reset counter
			phy_reset_counter <= 32'd0;
			
			// no reset performed yet
			phy_reset_performed <= 0;
			
			// assert the reset pin to trigger a reset of the PHY
			RST_reg <= 1;
			
			// do not register write while the PHY resets
			ulpi_register_write_reg <= 0;
			
			//led <= 4'b0000;
			//outdata <= 8'h8a;
		end
		
		//if (phy_reset_counter == 60000000)
		//if (phy_reset_counter == 10000000)
		if (phy_reset_counter == 1000000)
		begin
		
			
		
			phy_reset_counter <= 0;
			
			// YORO - you only reset once
			if (phy_reset_performed == 0)
			begin
`ifdef USE_LED_FOR_RESET_BLOCK
				led <= ~4'b1100;
`endif
			
				// PHY reset has been performed
				phy_reset_performed <= 1;
				
				// do not reset any more
				RST_reg <= 0;
				
				// start register write
				ulpi_register_write_reg <= 1;
				
			end
			
		end
		else
		begin
		
			phy_reset_counter <= phy_reset_counter + 32'd1;
			
		end		
		
	end
	
	
	
	
	
	
	
	
	
	//
	// Config State Machine 
	// - disables OTG activating peripheral mode
	// - enable Fast Speed (FS) mode by writing 0x45 into the FUNC_CTRL register
	//
	
	localparam CONFIG_STATE_0 		= 8'd0;
	localparam CONFIG_STATE_1 		= 8'd1;
	localparam CONFIG_STATE_2 		= 8'd2;
	localparam CONFIG_STATE_3 		= 8'd3;
	localparam CONFIG_STATE_4 		= 8'd4;
	localparam CONFIG_STATE_5 		= 8'd5;
	localparam CONFIG_STATE_6 		= 8'd6;
	localparam CONFIG_STATE_7 		= 8'd7;
	localparam CONFIG_STATE_8 		= 8'd8;
	localparam CONFIG_STATE_9 		= 8'd9;
	
	localparam CONFIG_STATE_10 	= 8'd10;
	localparam CONFIG_STATE_11		= 8'd11;
	localparam CONFIG_STATE_12		= 8'd12;
	localparam CONFIG_STATE_13		= 8'd13;
	localparam CONFIG_STATE_14		= 8'd14;
	localparam CONFIG_STATE_15		= 8'd15;
	localparam CONFIG_STATE_16		= 8'd16;	
	
	localparam MSG_DEV_DESC_0		= 8'd20;
	localparam MSG_DEV_DESC_1		= 8'd21;	
	localparam MSG_DEV_DESC_2		= 8'd22;	
	localparam MSG_DEV_DESC_3		= 8'd23;
	localparam MSG_DEV_DESC_4		= 8'd24;
	localparam MSG_DEV_DESC_5		= 8'd25;
	localparam MSG_DEV_DESC_6		= 8'd26;
	localparam MSG_DEV_DESC_7		= 8'd27;
	localparam MSG_DEV_DESC_8		= 8'd28;
	localparam MSG_DEV_DESC_9		= 8'd29;
	
	localparam MSG_DEV_DESC_10		= 8'd30;
	localparam MSG_DEV_DESC_11		= 8'd31;
	localparam MSG_DEV_DESC_12		= 8'd32;
	localparam MSG_DEV_DESC_13		= 8'd33;	
	localparam MSG_DEV_DESC_14		= 8'd34; // PID IN detection starts here
	localparam MSG_DEV_DESC_15		= 8'd35;
	localparam MSG_DEV_DESC_16		= 8'd36;
	localparam MSG_DEV_DESC_17		= 8'd37;
	localparam MSG_DEV_DESC_18		= 8'd38;
	localparam MSG_DEV_DESC_19		= 8'd39;
	
	localparam MSG_DEV_DESC_20		= 8'd40;
	localparam MSG_DEV_DESC_21		= 8'd41;
	localparam MSG_DEV_DESC_22		= 8'd42;
	localparam MSG_DEV_DESC_23		= 8'd43;
	localparam MSG_DEV_DESC_24		= 8'd44;
	localparam MSG_DEV_DESC_25		= 8'd45;
	localparam MSG_DEV_DESC_26		= 8'd46;
	localparam MSG_DEV_DESC_27		= 8'd47;
	localparam MSG_DEV_DESC_28		= 8'd48;
	localparam MSG_DEV_DESC_29		= 8'd49;
	
	localparam MSG_DEV_DESC_30		= 8'd50;
	localparam MSG_DEV_DESC_31		= 8'd51;
	localparam MSG_DEV_DESC_32		= 8'd52;
	localparam MSG_DEV_DESC_33		= 8'd53;
	localparam MSG_DEV_DESC_34		= 8'd54;
	localparam MSG_DEV_DESC_35		= 8'd55;
	localparam MSG_DEV_DESC_36		= 8'd56;
	localparam MSG_DEV_DESC_37		= 8'd57;
	localparam MSG_DEV_DESC_38		= 8'd58;
	localparam MSG_DEV_DESC_39		= 8'd59;
	
	localparam MSG_DEV_DESC_40		= 8'd60;
	localparam MSG_DEV_DESC_41		= 8'd61;
	localparam MSG_DEV_DESC_42		= 8'd62;
	localparam MSG_DEV_DESC_43		= 8'd63;
	localparam MSG_DEV_DESC_44		= 8'd64;
	localparam MSG_DEV_DESC_45		= 8'd65;
	localparam MSG_DEV_DESC_46		= 8'd66;
	localparam MSG_DEV_DESC_47		= 8'd67;
	localparam MSG_DEV_DESC_48		= 8'd68;
	localparam MSG_DEV_DESC_49		= 8'd69;
	
	localparam MSG_DEV_DESC_50		= 8'd70;
	localparam MSG_DEV_DESC_51		= 8'd71;
	localparam MSG_DEV_DESC_52		= 8'd72;
	localparam MSG_DEV_DESC_53		= 8'd73;
	localparam MSG_DEV_DESC_54		= 8'd74;
	localparam MSG_DEV_DESC_55		= 8'd75;
	localparam MSG_DEV_DESC_56		= 8'd76;
	localparam MSG_DEV_DESC_57		= 8'd77;
	localparam MSG_DEV_DESC_58		= 8'd78;
	localparam MSG_DEV_DESC_59		= 8'd79;
	
	localparam MSG_DEV_DESC_60		= 8'd80;
	localparam MSG_DEV_DESC_61		= 8'd81;
	localparam MSG_DEV_DESC_62		= 8'd82;
	localparam MSG_DEV_DESC_63		= 8'd83;
	localparam MSG_DEV_DESC_64		= 8'd84;
	localparam MSG_DEV_DESC_65		= 8'd85;
	localparam MSG_DEV_DESC_66		= 8'd86;
	localparam MSG_DEV_DESC_67		= 8'd87;
	localparam MSG_DEV_DESC_68		= 8'd88;
	localparam MSG_DEV_DESC_69		= 8'd89;
	
	localparam MSG_DEV_DESC_70		= 8'd90;
	localparam MSG_DEV_DESC_71		= 8'd91;
	localparam MSG_DEV_DESC_72		= 8'd92;
	localparam MSG_DEV_DESC_73		= 8'd93;
	localparam MSG_DEV_DESC_74		= 8'd94;
	localparam MSG_DEV_DESC_75		= 8'd95;
	localparam MSG_DEV_DESC_76		= 8'd96;
	localparam MSG_DEV_DESC_77		= 8'd97;
	localparam MSG_DEV_DESC_78		= 8'd98;
	localparam MSG_DEV_DESC_79		= 8'd99;
	
	localparam MSG_DEV_DESC_80		= 8'd100;
	localparam MSG_DEV_DESC_81		= 8'd101;
	localparam MSG_DEV_DESC_82		= 8'd102;
	localparam MSG_DEV_DESC_83		= 8'd103;
	localparam MSG_DEV_DESC_84		= 8'd104;
	localparam MSG_DEV_DESC_85		= 8'd105;
	localparam MSG_DEV_DESC_86		= 8'd106;
	localparam MSG_DEV_DESC_87		= 8'd107;
	localparam MSG_DEV_DESC_88		= 8'd108;
	localparam MSG_DEV_DESC_89		= 8'd109;
	
	localparam MSG_DEV_DESC_90		= 8'd110;
	localparam MSG_DEV_DESC_91		= 8'd111;
	localparam MSG_DEV_DESC_92		= 8'd112;
	localparam MSG_DEV_DESC_93		= 8'd113;
	localparam MSG_DEV_DESC_94		= 8'd114;
	localparam MSG_DEV_DESC_95		= 8'd115;
	localparam MSG_DEV_DESC_96		= 8'd116;
	localparam MSG_DEV_DESC_97		= 8'd117;
	localparam MSG_DEV_DESC_98		= 8'd118;
	localparam MSG_DEV_DESC_99		= 8'd119;
	
	localparam MSG_DEV_DESC_100		= 8'd120;
	localparam MSG_DEV_DESC_101		= 8'd121;
	localparam MSG_DEV_DESC_102		= 8'd122;
	localparam MSG_DEV_DESC_103		= 8'd123;
	localparam MSG_DEV_DESC_104		= 8'd124;
	localparam MSG_DEV_DESC_105		= 8'd125;
	localparam MSG_DEV_DESC_106		= 8'd126;
	localparam MSG_DEV_DESC_107		= 8'd127;
	localparam MSG_DEV_DESC_108		= 8'd128;
	localparam MSG_DEV_DESC_109		= 8'd129;
	
	localparam MSG_DEV_DESC_CENTER		= 8'hFE;
	
	localparam STATE_IDLE 			= 8'd255;
	
	reg [7:0] state;// <= STATE_IDLE;
	
	// combinational always block for next state logic
	//always @(config_cur_state)
	always @(posedge CLKOUT)	
	begin
	
		// default next state assignment
		//state = STATE_IDLE;
		
		if (!reset) 
		begin
			state = STATE_IDLE;
		end

		case (state)

			CONFIG_STATE_0: 
			begin			
`ifdef USE_LED_FOR_CONFIG_BLOCK
				//led_reg <= ~4'b0000;
				//led <= led_reg;
				led <= ~4'b0001;
`endif

				// LINK needs to pull STP low otherwise nothing works at all
				STP = 1'b0;

				if (DIR == 1)
				begin
					state <= CONFIG_STATE_0;
				end
				else
				begin

					// A ULPI READ is described by 11xxxxxx in binary. The xxxxxx contains the address. 
					// To read Vendor ID Low, the address is 0x00. So combining the CMD BITS with the address 
					// 0x00 yields 11000000b = 0xC0.
					// 11000000bin = 0xC0
					
					//outdata = 8'hC0; 	// vendor id low  	(0x24, 00100100) (ULPI register READ: address 0x00)
					//outdata = 8'hC1; 	// vendor id high 	(0x04, 00000100) (ULPI register READ: address 0x01)
					
					//outdata = 8'hC2; 		// product id low  	(0x04, 00000100) (ULPI register READ: address 0x02)
					//outdata = 8'hC3; 	// product id high 	(0x00, 00000000) (ULPI register READ: address 0x03)
					
					//outdata = 8'hC4; // function control
					
					//outdata = 8'hCD; // USB Interrupt Enable Rising
					
					//outdata = 8'hD3;
					
					// A ULPI WRITE 
					
					// https://cross-hair.co.uk/tech-articles/ULPI%20interface.html
					// First we must disable OTG features by writing x"00" to the OTG_CTRL (x"0a") register.
					// A TXCMD byte of x"8a" is sent then a data byte of x"00" as per Figure 1.
					
					outdata <= 8'h8a; // [10][0x0A]
					
					state <= CONFIG_STATE_1; // next state
				end
			end

			CONFIG_STATE_1:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b0001;
`endif
				outdata <= 8'h8a; // [10][0x0A]
				
				state <= CONFIG_STATE_2; // next state
			end
			
			CONFIG_STATE_2:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				//led_reg <= ~4'b0010;
				//led <= led_reg;
				led <= ~4'b0010;
`endif
				// write to the OTG register
				outdata <= 8'h8a; // [10][0x0A]
				
				state <= CONFIG_STATE_3; // next state
			end
			
			CONFIG_STATE_3:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				//led_reg <= ~4'b0011;
				//led <= led_reg;
				led <= ~4'b0011;
`endif
				outdata <= 8'h00; // data byte to write into the register
				
				state <= CONFIG_STATE_4; // next state
			end
			
			CONFIG_STATE_4:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				//led_reg <= ~4'b0100;
				//led <= led_reg;
				led <= ~4'b0100;
`endif
				// write 0x00 to the OTG register to disable OTG and enable peripheral mode
				outdata <= 8'h00;
				STP <= 1'b1; // send STP to tell the PHY that the command is sent completely and no more bytes follow
			
				state <= CONFIG_STATE_5; // next state
			end
			
			CONFIG_STATE_5:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK	
				//led_reg <= ~4'b0101;
				//led <= led_reg;
				led <= ~4'b0101;
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
			
				state <= CONFIG_STATE_6; // next state
			end
			
			CONFIG_STATE_6:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b0110;
`endif
				// Write to the FUNC_CTRL register (Goal: enable Fast Speed (FS) mode)
				outdata <= 8'h84; // [10][0x04] write the function control register
					
				state <= CONFIG_STATE_7; // next state
			end 
			
			CONFIG_STATE_7:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b0110;
`endif
				// Write to the FUNC_CTRL register (Goal: enable Fast Speed (FS) mode)
				outdata <= 8'h84; // [10][0x04] write the function control register
					
				state <= CONFIG_STATE_8; // next state
			end
			
			CONFIG_STATE_8:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b1000;
`endif
				// Write to the FUNC_CTRL register (Goal: enable Fast Speed (FS) mode)
				outdata <= 8'h84; // [10][0x04] write the function control register
					
				state <= CONFIG_STATE_9; // next state
			end
			
			CONFIG_STATE_9:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b0000;
`endif
				// write the value 0x45 into the FUNC_CTRL register to enable Fast Speed (FS) mode.
				outdata <= 8'h45; // data byte to write into the register (0100 0101)
					
				state <= CONFIG_STATE_10; // next state
			end
			
			CONFIG_STATE_10:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b1010;
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
				
				// The PHY should respond with a RXCMD showing a LineState of J ("01", FS Idle).
				// 10001010
					
				state <= CONFIG_STATE_11; // next state
			end
			
			CONFIG_STATE_11:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b0011;
`endif
				outdata <= 8'h00;
				STP <= 1'b1; // send STP to tell the PHY that the command is sent completely and no more bytes follow
					
				state <= CONFIG_STATE_12; // next state
			end
			
			CONFIG_STATE_12:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b1100;
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
					
				state <= CONFIG_STATE_13; // next state
			end
			
			CONFIG_STATE_13:
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b1101;
`endif
				//outdata = 8'b01000000; // Transmit on D+/D- (See Table 6.4, page 24) [01]
				//STP = 8'h00;
				
				outdata <= 8'h00;
				STP <= 1'b0;
				
				state <= CONFIG_STATE_14; // next state
			end
			
			CONFIG_STATE_14:
			begin			
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b1110;
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
					
				state <= MSG_DEV_DESC_0;		
			end
			
			
			
			CONFIG_STATE_16:
			begin
				state <= CONFIG_STATE_16;
			end
			
			
			
			//default:
			//begin				
				// next state
			//	state <= CONFIG_IDLE; // Fallback to default state
				
				// LINK needs to pull STP low otherwise nothing works at all
			//	STP <= 0;
			//end			
			
		//endcase

	//end	
	
	//always @(posedge CLKOUT)
	//begin
	
		//if (!reset)
		//begin
		//	state = MSG_DEV_DESC_0;
		//end
	
		//case (state)
		
		
		
			MSG_DEV_DESC_CENTER:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1101;
`endif
				if (data == 8'hC3) // 0xC3 is 1100 0011 == PID DATA 0
					// CONSUME: GetDescriptor
					state <= MSG_DEV_DESC_1;
				//else if (data == 8'hE1)
					// CONSUME: PID OUT <E1 00 10> (Send after RESPONSE to GetDescriptor, 
				//	state <= MSG_DEV_DESC_41;
				//else if (data == 8'hC3)	// PID DATA0 - 0xC3 11000011 // mystery packet
				//	state <= MSG_DEV_DESC_50;
				//else if (data == 8'h4B)
				//	state <= MSG_DEV_DESC_44;
				else
					state <= MSG_DEV_DESC_CENTER;
			end
			
			
			//
			// SET ADDRESS 00 05 (03|04) 00 00 00 00 00
			// 
			
			MSG_DEV_DESC_90:
			begin
				if (data == 8'h05)
				begin
					state <= MSG_DEV_DESC_91;
				end
				else
					state <= MSG_DEV_DESC_90;
			end
			
			MSG_DEV_DESC_91:
			begin
				if (data == 8'h03)
				begin
					state <= MSG_DEV_DESC_92;
				end
				else if (data == 8'h04)
				begin
					state <= MSG_DEV_DESC_92;
				end
				else
					state <= MSG_DEV_DESC_91;
			end
			
			MSG_DEV_DESC_92:
			begin
				if (data == 8'h00)
				begin
					state <= MSG_DEV_DESC_93;
				end
				else
					state <= MSG_DEV_DESC_92;
			end
			
			MSG_DEV_DESC_93:
			begin
				if (data == 8'h00)
				begin
					state <= MSG_DEV_DESC_94;
				end
				else
					state <= MSG_DEV_DESC_93;
			end
			
			MSG_DEV_DESC_94:
			begin
				if (data == 8'h00)
				begin
					state <= MSG_DEV_DESC_95;
				end
				else
					state <= MSG_DEV_DESC_94;
			end
			
			MSG_DEV_DESC_95:
			begin
				if (data == 8'h00)
				begin
					state <= MSG_DEV_DESC_96;
				end
				else
					state <= MSG_DEV_DESC_95;
			end
			
			MSG_DEV_DESC_96:
			begin
				if (data == 8'h00)
				begin
					state <= MSG_DEV_DESC_97;
				end
				else
					state <= MSG_DEV_DESC_96;
			end
			
			// CRC 1
			MSG_DEV_DESC_97:
			begin
				state <= MSG_DEV_DESC_98;
			end
			
			// CRC 2
			MSG_DEV_DESC_98:
			begin
				state <= MSG_DEV_DESC_99;
			end
			
			//
			// SEND ACK
			//
			// Wait for the PHY to release the lines and send ACK (0x42)
			// The PHY will produce the SYNC pattern and the EOP for us!!! THANK YOU!
			//
			
			MSG_DEV_DESC_99:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0011; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_99;
				end
				else 
				begin
					outdata <= 8'h42; // ack 0x42 == [01] 00 0010
					STP <= 1'b0;
					
					state <= MSG_DEV_DESC_100;
				end				
			end
			
			MSG_DEV_DESC_100:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1100; // [L1][L2][L3][L4]
`endif
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_100;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b1;
						state <= MSG_DEV_DESC_101;
					end
					else 
						state <= state;
			end
			
			MSG_DEV_DESC_101:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1101; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
				state <= MSG_DEV_DESC_102;
				//state <= MSG_DEV_DESC_CENTER;
			end
			
			//
			// CONSUME PID IN 69
			//
			
			MSG_DEV_DESC_102:
			begin
				if (data == 8'h69)
				begin
					state <= MSG_DEV_DESC_103;
				end
				else
					state <= MSG_DEV_DESC_102;
			end
			
			// ADDR ENDP
			MSG_DEV_DESC_103:
			begin
				state <= MSG_DEV_DESC_104;
			end
			
			// CRC6
			MSG_DEV_DESC_104:
			begin
				state <= MSG_DEV_DESC_105;
			end
			
			//
			// SEND DATA 1 [4B 00 00]
			//
		
			MSG_DEV_DESC_105:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0011; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_105;
				end
				else 
				begin
					outdata <= 8'h4B; // ack 0x4B == [01] 00 1001
					STP <= 1'b0;
					
					state <= MSG_DEV_DESC_106;
				end				
			end
			
			MSG_DEV_DESC_106:
			begin
				if (DIR == 1)
					state <= MSG_DEV_DESC_106;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b0;
						state <= MSG_DEV_DESC_107;
					end
					else 
						state <= state;
			end
			
			MSG_DEV_DESC_107:
			begin
				if (DIR == 1)
					state <= MSG_DEV_DESC_107;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b0;
						state <= MSG_DEV_DESC_108;
					end
					else 
						state <= state;
			end
			
			MSG_DEV_DESC_108:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1100; // [L1][L2][L3][L4]
`endif
/**/
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_108;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b1;
						state <= MSG_DEV_DESC_109;
					end
					else 
						state <= state;

//				// tell the phy that the outgoing message is completely output
//				outdata <= 8'h00;
//				STP <= 1'b1;
//				state <= MSG_DEV_DESC_109;
			end
			
			MSG_DEV_DESC_109:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1101; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
				//state <= MSG_DEV_DESC_102;
				state <= MSG_DEV_DESC_CENTER;
			end
			
			//
			// CONSUME GET_DESCRIPTOR_REQUEST
			// 80 06 00 01 00 00 40 00
			//
			// CONSUME SET_ADDRESS
			// 00 05 03 00 00 00 00 00 <
			// 
			
			MSG_DEV_DESC_1:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001;
`endif
//				if (data == 8'h80) // [80] 
//					state <= MSG_DEV_DESC_2;
//				else if (data == 8'h00) // [00] 05 03 00 00 00 00 00
//					state <= MSG_DEV_DESC_90;
//				else
//					state <= MSG_DEV_DESC_1;
					
				case (data)
				
					8'h80:
					begin
						state <= MSG_DEV_DESC_2;
					end
					
					8'h00:
					begin
						state <= MSG_DEV_DESC_90;
					end
					
					default:
					begin
						state <= MSG_DEV_DESC_1;
					end
					
				endcase
				
			end
			
			MSG_DEV_DESC_2:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0010;
`endif
				if (data == 8'h06) // <80 [06]
					state <= MSG_DEV_DESC_3;
				else
					state <= MSG_DEV_DESC_2;
			end
			
			MSG_DEV_DESC_3:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0011; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// <80 06 [00]
					state <= MSG_DEV_DESC_4;
				else
					state <= MSG_DEV_DESC_3;
			end
			
			MSG_DEV_DESC_4:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0100; // [L1][L2][L3][L4]
`endif
				if (data == 8'h01)  // <80 06 00 [01]
					state <= MSG_DEV_DESC_5;
				else
					state <= MSG_DEV_DESC_4;
			end
			
			MSG_DEV_DESC_5:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0101; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// <80 06 00 01 [00]
					state <= MSG_DEV_DESC_6;
				else
					state <= MSG_DEV_DESC_5;
			end
			
			MSG_DEV_DESC_6:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0110; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// <80 06 00 01 00 [00]
					state <= MSG_DEV_DESC_7;
				else
					state <= MSG_DEV_DESC_6;
			end
			
			MSG_DEV_DESC_7:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0110; // [L1][L2][L3][L4]
`endif
				if (data == 8'h40)	// <80 06 00 01 00 00 [40]
					state <= MSG_DEV_DESC_8;
				else if (data == 8'h12)
					state <= MSG_DEV_DESC_8;
				else
					state <= MSG_DEV_DESC_7;
			end
			
			MSG_DEV_DESC_8:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1000; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// <80 06 00 01 00 00 40 [00]> <DD 94>
					state <= MSG_DEV_DESC_9; // entire DEVICE DESCRIPTOR REQUEST PACKET RECEIVED
				else
					state <= MSG_DEV_DESC_8;
			end
			
			//
			// CRC16 (2 Byte CRC) which we consume but skip checking validity
			//
			
			MSG_DEV_DESC_9:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif
				state <= MSG_DEV_DESC_10; // SKIP CRC BYTE 0
			end
			
			MSG_DEV_DESC_10:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1010; // [L1][L2][L3][L4]
`endif
				state <= MSG_DEV_DESC_11; // SKIP CRC BYTE 1
			end
			
			//
			// SEND ACK
			//
			// Wait for the PHY to release the lines and send ACK (0x42)
			// The PHY will produce the SYNC pattern and the EOP for us!!! THANK YOU!
			//
			
			MSG_DEV_DESC_11:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0011; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_11;
				end
				else 
				begin
					outdata <= 8'h42; // ack 0x42 == [01] 00 0010
					STP <= 1'b0;
					
					state <= MSG_DEV_DESC_12;
				end
				
			end
			
			MSG_DEV_DESC_12:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1100; // [L1][L2][L3][L4]
`endif
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_12;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b1;
						state <= MSG_DEV_DESC_13;
					end
				else 
					state <= state;
			end
			
			MSG_DEV_DESC_13:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1101; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
				state <= MSG_DEV_DESC_14;
			end
			
			//
			// CONSUME PID IN
			//
			// PID IN detection starts here. We expect the bytes <BYTES: 69 00 10>
			//
			
			MSG_DEV_DESC_14:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1110; // [L1][L2][L3][L4]
`endif
				if (data == 8'h69) // PID BYTE 0 - 0x69
					state <= MSG_DEV_DESC_15;
				else
					state <= MSG_DEV_DESC_14;
			end
			
			MSG_DEV_DESC_15:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1110; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 1 - 0x00
					state <= MSG_DEV_DESC_16;
				else
					state <= MSG_DEV_DESC_15;
			end
			
			MSG_DEV_DESC_16:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1110; // [L1][L2][L3][L4]
`endif
				if (data == 8'h10)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_17;
				else
					state <= MSG_DEV_DESC_16;
			end
			
			//
			// SEND device descriptor
			//
			
			MSG_DEV_DESC_17:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_17; // remain
				end
				else 
				begin
					// 0x4B == 01 00 1011
					outdata <= 8'h4B; // <[4B] 12 01 00 02 FF FF FF 40 DE AD BE EF 01 00 00 00 00 01>
					STP <= 1'b0;					
					state <= MSG_DEV_DESC_18; // next state
				end		
			end
			MSG_DEV_DESC_18:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_18; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// length of descriptor
						outdata <= 8'h12; // <4B [12] 01 00 02 FF FF FF 40 DE AD BE EF 01 00 00 00 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_19; // next state
					end
					else 
						state <= state;
				end				
			end
			MSG_DEV_DESC_19:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_19; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// descriptor type 
						outdata <= 8'h01; // <4B 12 [01] 00 02 FF FF FF 40 DE AD BE EF 01 00 00 00 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_20; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_20:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_20; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// usb version
						//outdata <= 8'h00; // <4B 12 01 [00] 02 FF FF FF 40 DE AD BE EF 01 00 00 00 00 01>
						outdata <= 8'h10;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_21; // next state
					end
					else 
						state <= state;
				end						
			end
			MSG_DEV_DESC_21:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_21; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// usb version
						
						//outdata <= 8'h02; // <4B 12 01 00 [02] FF FF FF 40 DE AD BE EF 01 00 00 00 00 01>
						outdata <= 8'h01;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_22; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_22:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_22; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// device Class
						
						//outdata <= 8'hFF; // <4B 12 01 00 02 [FF] FF FF 40 DE AD BE EF 01 00 00 00 00 01>
						outdata <= 8'h00; 
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_23; // next state
					end
					else 
						state <= state;
				end				
			end
			MSG_DEV_DESC_23:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_23; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// device subclass
						
						//outdata <= 8'hFF; // <4B 12 01 00 02 FF [FF] FF 40 DE AD BE EF 01 00 00 00 00 01>
						outdata <= 8'h00;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_24; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_24:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// Wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_24; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// device protocol
						//outdata <= 8'hFF; // <4B 12 01 00 02 FF FF [FF] 40 DE AD BE EF 01 00 00 00 00 01>
						outdata <= 8'h00;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_25; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_25:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_25; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// bMaxPacketSize0 == 8 (8 bytes)
						outdata <= 8'h40; // <4B 12 01 00 02 FF FF FF [40] DE AD BE EF 01 00 00 00 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_26; // next state
					end
					else 
						state <= state;
				end					
			end			
			MSG_DEV_DESC_26:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif	
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_26; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// id vendor 1
						//outdata <= 8'hDE; // <4B 12 01 00 02 FF FF FF 40 [DE] AD BE EF 01 00 00 00 00 01>
						outdata <= 8'hC4;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_27; // next state
					end
					else 
						state <= state;
				end			
			end			
			MSG_DEV_DESC_27:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_27; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// id vendor 2
						//outdata <= 8'hAD; // <4B 12 01 00 02 FF FF FF 40 DE [AD] BE EF 01 00 00 00 00 01>
						outdata <= 8'h10; 
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_28; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_28:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_28; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// id product 1
						//outdata <= 8'hBE; // <4B 12 01 00 02 FF FF FF 40 DE AD [BE] EF 01 00 00 00 00 01>
						outdata <= 8'h60;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_29; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_29:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_29; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// id product 2
						//outdata <= 8'hEF; // <4B 12 01 00 02 FF FF FF 40 DE AD BE [EF] 01 00 00 00 00 01>
						outdata <= 8'hEA;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_30; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_30:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_30; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// bcdDevice (1/2)
						outdata <= 8'h00; // <4B 12 01 00 02 FF FF FF 40 DE AD BE EF [01] 00 00 00 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_31; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_31:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_31; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// bcdDevice (2/2)
						outdata <= 8'h01; // <4B 12 01 00 02 FF FF FF 40 DE AD BE EF 01 [00] 00 00 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_32; // next state
					end
					else 
						state <= state;
				end					
			end			
			MSG_DEV_DESC_32:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_32; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// string descriptor 1
						outdata <= 8'h00; // <4B 12 01 00 02 FF FF FF 40 DE AD BE EF 01 00 [00] 00 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_33; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_33:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_33; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// string descriptor 2
						outdata <= 8'h00; // <4B 12 01 00 02 FF FF FF 40 DE AD BE EF 01 00 00 [00] 00 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_34; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_34:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_34; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// string descriptor 3
						outdata <= 8'h00; // <4B 12 01 00 02 FF FF FF 40 DE AD BE EF 01 00 00 00 [00] 01>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_35; // next state
					end
					else 
						state <= state;
				end					
			end
			MSG_DEV_DESC_35:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_35; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// bNumConfigurations
						outdata <= 8'h01; // <4B 12 01 00 02 FF FF FF 40 DE AD BE EF 01 00 00 00 00 [01]>
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_36; // next state
					end
					else 
						state <= state;
				end					
			end			
			MSG_DEV_DESC_36:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_36; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// CRC 1
						//outdata <= 8'hC0; // <4B 12 01 00 02 FF FF FF 08 33 16> THE CRC IS PROVIDED IN REVERSE!!!! 16 first
						outdata <= 8'hDB;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_37; // next state
					end
					else 
						state <= state;
				end
			end
			MSG_DEV_DESC_37:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif			
				// wait for the line to be free
				if (DIR == 1)
				begin
					state <= MSG_DEV_DESC_37; // remain
				end
				else 
				begin
					if (NXT == 1)
					begin
						// CRC 2
						//outdata <= 8'hCE; // <4B 12 01 00 02 FF FF FF 08 33 16> THE CRC IS PROVIDED IN REVERSE!!!! 33 last
						outdata <= 8'h34;
						STP <= 1'b0;					
						state <= MSG_DEV_DESC_38; // next state
					end
					else 
						state <= state;
				end			
			end
			
			// SET STOP BIT
			MSG_DEV_DESC_38:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1100; // [L1][L2][L3][L4]
`endif
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_38;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b1;						
						state <= MSG_DEV_DESC_39;
					end
					else 
						state <= MSG_DEV_DESC_38;

//				// tell the phy that the outgoing message is completely output
//				outdata <= 8'h00;
//				STP <= 1'b1;						
//				state <= MSG_DEV_DESC_39;
			end
			
			// REMOVE the stop bit
			MSG_DEV_DESC_39:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0110; // [L1][L2][L3][L4]
`endif		
				outdata <= 8'h00;
				STP <= 1'b0;
				state <= MSG_DEV_DESC_40;
			end
			
			
			
			
			
			// CONSUME ACK
			MSG_DEV_DESC_40:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0000; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
				if (data == 8'hD2)
					state <= MSG_DEV_DESC_41;
				else
					state <= MSG_DEV_DESC_40;
			end
			
			
			
			
			
			
			//
			// CONSUME: PID OUT <E1 00 10>
			//

			MSG_DEV_DESC_41:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0000; // [L1][L2][L3][L4]
`endif
				if (data == 8'hE1) // PID BYTE 0
					state <= MSG_DEV_DESC_42;
				else
					state <= MSG_DEV_DESC_41;
			end

			MSG_DEV_DESC_42:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0001; // [L1][L2][L3][L4]
`endif
				//if (data == 8'h00)	// PID BYTE 1 - 0x00
				//	state <= MSG_DEV_DESC_43;
				//else
				//	state <= MSG_DEV_DESC_42;
				state <= MSG_DEV_DESC_43;
			end
			
			MSG_DEV_DESC_43:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0010; // [L1][L2][L3][L4]
`endif
				//if (data == 8'h10)	// PID BYTE 2 - 0x10
				//	state <= MSG_DEV_DESC_44;
				//else
				//	state <= MSG_DEV_DESC_43;
				state <= MSG_DEV_DESC_44;
			end
			
			//
			// CONSUME: PID DATA 1 <4B 00 00>
			//
			
			MSG_DEV_DESC_44:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0100; // [L1][L2][L3][L4]
`endif
				if (data == 8'h4D) // PID BYTE 0 - 0x4B [01][00][1011]
					state <= MSG_DEV_DESC_45;
				//if (data == 8'h4B) // PID BYTE 0 - 0x4B [01][00][1011]
				//	state <= MSG_DEV_DESC_44;
				else
					state <= MSG_DEV_DESC_44;
			end
			
			MSG_DEV_DESC_45:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0101; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 1 - 0x00
					state <= MSG_DEV_DESC_46;
				else
					state <= MSG_DEV_DESC_45;
			end
			
			MSG_DEV_DESC_46:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0110; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x00
					state <= MSG_DEV_DESC_47;
				else
					state <= MSG_DEV_DESC_46;
			end
			
			//
			// SEND: ACK <D2>
			//
			// Wait for the PHY to release the lines and send ACK (0x42)
			// The PHY will produce the SYNC pattern and the EOP for us!!! THANK YOU!
			//
			
			MSG_DEV_DESC_47:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1010; // [L1][L2][L3][L4]
`endif		
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_47;
				end
				else 
				begin
					outdata <= 8'h42; // ack (01000010)
					STP <= 1'b0;
					
					state <= MSG_DEV_DESC_48;
				end
			
			end
			
			MSG_DEV_DESC_48:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1000; // [L1][L2][L3][L4]
`endif
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_48;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						outdata <= 8'h00;
						STP <= 1'b1;
						state <= MSG_DEV_DESC_49;
					end
					else 
						state <= MSG_DEV_DESC_48;
			end
			
			// REMOVE the stop bit
			MSG_DEV_DESC_49:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1001; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0;
				
				//state <= MSG_DEV_DESC_49;
				state <= MSG_DEV_DESC_CENTER;
				
			end
			
			//
			// process the mystery request that the internet does not know ???
			// [PID DATA 0: C3] [00 05 03 00 00 00 00 00] [CRC: C7EA]
			//
			
			MSG_DEV_DESC_49:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1000; // [L1][L2][L3][L4]
`endif
				if (data == 8'hC3)	// PID DATA 0 - 0xC3 11000011
					state <= MSG_DEV_DESC_50;
				else
					state <= MSG_DEV_DESC_49;
			end
			
			MSG_DEV_DESC_50:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1001; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_51;
				else
					state <= MSG_DEV_DESC_50;
			end
			MSG_DEV_DESC_51:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1001; // [L1][L2][L3][L4]
`endif
				if (data == 8'h05)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_52;
				else
					state <= MSG_DEV_DESC_51;
			end
			MSG_DEV_DESC_52:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0000; // [L1][L2][L3][L4]
`endif
				if (data == 8'h03)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_53;
				else
					state <= MSG_DEV_DESC_52;
			end
			MSG_DEV_DESC_53:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0011; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_54;
				else
					state <= MSG_DEV_DESC_53;
			end
			MSG_DEV_DESC_54:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0100; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_55;
				else
					state <= MSG_DEV_DESC_54;
			end
			MSG_DEV_DESC_55:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0101; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_56;
				else
					state <= MSG_DEV_DESC_55;
			end
			MSG_DEV_DESC_56:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0000; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_57;
				else
					state <= MSG_DEV_DESC_56;
			end
			MSG_DEV_DESC_57:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0101; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_58;
				else
					state <= MSG_DEV_DESC_57;
			end
			
			//
			// Consume CRC
			//
/*
			MSG_DEV_DESC_47:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0111; // [L1][L2][L3][L4]
`endif
				if (data == 8'hEA)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_48;
				else
					state <= MSG_DEV_DESC_47;
			end
			MSG_DEV_DESC_48:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0111; // [L1][L2][L3][L4]
`endif
				if (data == 8'hC7)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_49;
				else
					state <= MSG_DEV_DESC_48;
			end
*/

			//
			// CRC16 (2 Byte CRC) which we consume but skip checking validity
			//
			
			MSG_DEV_DESC_58:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1001; // [L1][L2][L3][L4]
`endif
				state <= MSG_DEV_DESC_59; // SKIP CRC BYTE 0
			end
			
			MSG_DEV_DESC_59:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1010; // [L1][L2][L3][L4]
`endif
				state <= MSG_DEV_DESC_60; // SKIP CRC BYTE 1
			end
			
			//
			// SEND ACK
			//
			// Wait for the PHY to release the lines and send ACK (0x42)
			// The PHY will produce the SYNC pattern and the EOP for us!!! THANK YOU!
			//
			
			MSG_DEV_DESC_60:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0111; // [L1][L2][L3][L4]
`endif		


				outdata <= 8'h42; // ack (READ: 6.1.7.6 Typical USB Transmit with ULPI in document: 00001783C.pdf)
				// a transmit command looks like this: [01][00][xxxx] whereas xxxx = 4 bit PID. The PID for
				// an acknowledge ACK is: 0010
				
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_60;
				end
				else 
				begin					
					STP <= 1'b0;					
					state <= MSG_DEV_DESC_61;
				end
			end
			
			MSG_DEV_DESC_61:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1000; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_61;
				else 
					if (NXT == 1)
					begin
						// tell the phy that the outgoing message is completely output
						STP <= 1'b1;
						state <= MSG_DEV_DESC_62;
					end
					else 
						state <= state;
			end
			
			// PULL STOP LOW
			MSG_DEV_DESC_62:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1011; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0; // pull the STP signal low because it is high for a single cycle only
				state <= MSG_DEV_DESC_63;
			end
			
			//
			// CONSUME: (Host -> Device) PID IN <69 00 10>
			//
			
			MSG_DEV_DESC_63:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1001; // [L1][L2][L3][L4]
`endif
				if (data == 8'h69) // PID BYTE 0 - 0x69
					state <= MSG_DEV_DESC_64;
				else
					state <= MSG_DEV_DESC_63;
			end
			
			MSG_DEV_DESC_64:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0000; // [L1][L2][L3][L4]
`endif
				if (data == 8'h00)	// PID BYTE 1 - 0x00
					state <= MSG_DEV_DESC_65;
				else
					state <= MSG_DEV_DESC_64;
			end
			
			MSG_DEV_DESC_65:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b0100; // [L1][L2][L3][L4]
`endif
				if (data == 8'h10)	// PID BYTE 2 - 0x10
					state <= MSG_DEV_DESC_66;
				else
					state <= MSG_DEV_DESC_65;
			end
			
			//
			// SEND: PID DATA 1 <00 00>
			//
			// Wait for the PHY to release the lines and send 0x00 0x00
			// The PHY will produce the SYNC pattern and the EOP for us!!! THANK YOU!
			//
			
			MSG_DEV_DESC_66:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1000; // [L1][L2][L3][L4]
`endif		

				//outdata <= 8'hD2; // ack 11 01 0010
				outdata <= 8'h4B; // ack (READ: 6.1.7.6 Typical USB Transmit with ULPI in document: 00001783C.pdf)
				// a transmit command looks like this: [01][00][xxxx] whereas xxxx = 4 bit PID. The PID for
				// an DATA 1 is: 1011
				//outdata <= 8'h4D; // ERROR Packet
				//outdata <= 8'h44;
				
				// Wait for the line to be free
				if (DIR || NXT)
				begin
					state <= MSG_DEV_DESC_66;
				end
				else 
				begin				
					STP <= 1'b0;					
					state <= MSG_DEV_DESC_67;
				end
			end
			
			MSG_DEV_DESC_67:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1001; // [L1][L2][L3][L4]
`endif		
				// WAIT for the DIR to be low so the line is not used
				if (DIR == 1)
					state <= MSG_DEV_DESC_67;
				else 
					if (NXT == 1)
					begin
						outdata <= 8'h00;
						// tell the phy that the outgoing message is completely output
						STP <= 1'b0;
						state <= MSG_DEV_DESC_68;
					end
					else 
						state <= state;
			end
			
			// PULL STOP LOW
			MSG_DEV_DESC_68:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1010; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 8'h00; // pull the STP signal low because it is high for a single cycle only
				state <= MSG_DEV_DESC_69;
			end
			
			// PULL STOP HIGH
			MSG_DEV_DESC_69:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1010; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b1; // pull the STP signal high because it is high for a single cycle only
				state <= MSG_DEV_DESC_70;
			end
			
			// PULL STOP LOW
			MSG_DEV_DESC_70:
			begin
`ifdef USE_LED_FOR_COMM_BLOCK
				led <= ~4'b1010; // [L1][L2][L3][L4]
`endif
				outdata <= 8'h00;
				STP <= 1'b0; // pull the STP signal low because it is high for a single cycle only
				state <= MSG_DEV_DESC_70;
			end
			
			STATE_IDLE: 
			begin
`ifdef USE_LED_FOR_CONFIG_BLOCK
				led <= ~4'b1000;
`endif
				// LINK needs to pull STP low otherwise nothing works at all
				STP <= 1'b0;
				
				// next state
				//if (ulpi_register_write_reg == 1)
				//begin
					//state <= CONFIG_STATE_0;
					state <= MSG_DEV_DESC_CENTER;
				//end
			end
			
			default:
				state <= STATE_IDLE;
			
		endcase
		
	end
	
endmodule